`timescale 1ns/1ps

module imem #(
    parameter int    XLEN        = riscv_pkg::XLEN,
    parameter int    DEPTH_WORDS = 64,
    parameter string MEMFILE     = ""          // optional: $readmemh file
    )(
    input  logic [XLEN-1:0] addr,              // byte address (PC)
    output logic [31:0]     r_d                // 32-bit instruction
    );
    import riscv_pkg::*;

    // ROM storage
    logic [31:0] mem [0:DEPTH_WORDS-1]; //fill addresses in increasing order

    // Optional preload from file; otherwise, hardcode
    initial begin
        // default NOPs to avoid Xs in sim
        for (int i = 0; i < DEPTH_WORDS; i++) mem[i] = INSTR_NOP;

        if (MEMFILE != "") begin
        $readmemh(MEMFILE, mem);
        end 
        else begin
        mem[0]  = 32'h0050_0113;
        mem[1]  = 32'h00C0_0193;
        mem[2]  = 32'hFF71_8393;
        mem[3]  = 32'h0023_E233;
        mem[4]  = 32'h0041_F2B3;
        mem[5]  = 32'h0042_82B3;
        mem[6]  = 32'h0272_8863;
        mem[7]  = 32'h0041_A233;
        mem[8]  = 32'h0002_0463;
        mem[9]  = 32'h0000_0293;
        mem[10] = 32'h0023_A233;
        mem[11] = 32'h0052_03B3;
        mem[12] = 32'h4023_83B3;
        mem[13] = 32'h0471_AA23;
        mem[14] = 32'h0600_2103;
        mem[15] = 32'h0051_04B3;
        mem[16] = 32'h0080_01EF;
        mem[17] = 32'h0010_0113;
        mem[18] = 32'h0091_0133;
        mem[19] = 32'h0221_A023;
        mem[20] = 32'h0021_0063;
        end
    end

    // Combinational ROM read
    assign r_d = mem[addr[31:2]];
endmodule
